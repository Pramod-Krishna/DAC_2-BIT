* /home/pramod/Desktop/esim/eSim-1.1.3/src/SubcircuitLibrary/r22/r22.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Aug  8 21:37:19 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad1_ eSim_MOS_P		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N		
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_M3-Pad3_ Net-_M3-Pad1_ eSim_MOS_P		
M4  Net-_M3-Pad3_ Net-_M1-Pad1_ Net-_M4-Pad3_ Net-_M4-Pad3_ eSim_MOS_N		
M6  Net-_M3-Pad3_ Net-_M1-Pad2_ Net-_M4-Pad3_ Net-_M3-Pad3_ eSim_MOS_P		
M5  Net-_M3-Pad1_ Net-_M1-Pad2_ Net-_M3-Pad3_ Net-_M3-Pad3_ eSim_MOS_N		
U1  Net-_M1-Pad2_ Net-_M4-Pad3_ Net-_M3-Pad1_ Net-_M3-Pad3_ PORT		
v1  Net-_M2-Pad1_ GND 3.3v		

.end
